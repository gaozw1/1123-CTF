    Mac OS X            	   2  �     �                                    ATTR;���  �   �   ?                  �   ?  com.apple.quarantine 0083;5bc985e7;DrUnarchiver;DFA483C0-F16F-479F-A025-FD1AD0310BF7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        This resource fork intentionally left blank                                                                                                                                                                                                                            ��